RLC LPF underdamped
*signal sources*
Vin 1 0 AC 1 0
*circuit description*
R1 1 2 10
L1 2 3 1000u
C1 3 0 100n
*AC analysis*
.AC DEC 200 1Hz 150kHz
* Output request
.PRINT AC V(1) V(3)
.PLOT AC V(1) V(3)



.end
