Linear Circuit


R1 1 2 20
 
R2 2 3 90

R3 3 4 80

R4 2 0 10

R6 3 0 40

Vb 1 0 40

Is 0 4 1

.op

.End
